* C:\Users\Mark\Documents\H-Bridge\H-Bridge.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/06/2016 2:16:27 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad3_ Net-_Q3-Pad3_ IRF540N		
Q6  Net-_Q5-Pad1_ Net-_Q5-Pad3_ Net-_Q3-Pad3_ IRF540N		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ IRF9540N		
Q5  Net-_Q5-Pad1_ Net-_Q2-Pad2_ Net-_Q5-Pad3_ IRF9540N		
R5  Net-_Q5-Pad3_ Net-_Q2-Pad3_ R		
Q4  Net-_Q4-Pad1_ Net-_Q3-Pad3_ GND IRF540N		
R4  Net-_Q4-Pad1_ ? 1M		
R2  Net-_Q2-Pad2_ Net-_Q1-Pad1_ 10k		
Q7  Net-_Q7-Pad1_ Net-_Q7-Pad2_ GND BC547		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ GND BC547		
R3  Net-_Q2-Pad1_ Net-_Q1-Pad1_ 1M		
R6  Net-_Q7-Pad1_ Net-_Q5-Pad1_ 1M		
R7  Net-_Q7-Pad1_ Net-_Q2-Pad2_ 10k		
R1  Net-_Q1-Pad2_ ? R		
R8  ? Net-_Q7-Pad2_ R		

.end
